-----------------------------------------------------------------------------------------------------------------------
-- Author:          Yu-Cheng Chen, ychen414@gatech.edu
--
-- Create Date:     16:43:30 09/02/2019
-- Module Name:     des_cipher_top_tb.vhd
-- Project Name:    des_cipher
-- Description:
--
--      Testbench for the des_cipher_top engine.
--      This is the testbench for the des_cipher_top engine. It exercises all the input control signals and error generation,
--      and tests the des_cipher_top engine.
--
-- Copyright: Georgia Institute of Technology 2019
--
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
--
--  Project structure:
--
--  |- des_cipher_top.vhd
--    |- des_top.vhd
--      |- block_top.vhd
--        |- add_key.vhd
--        |
--        |- add_left.vhd
--        |
--        |- e_expansion_function.vhd
--        |
--        |- p_box.vhd
--        |
--        |- s_box.vhd
--            |- s1_box.vhd
--            |- s2_box.vhd
--            |- s3_box.vhd
--            |- s4_box.vhd
--            |- s5_box.vhd
--            |- s6_box.vhd
--            |- s7_box.vhd
--            |- s8_box.vhd
--    |- key_schedule.vhd
-----------------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity des_cipher_top_tb is
    Generic (
        CLK_PERIOD : time := 10 ns                     -- clock period (default 100MHz)
    );
end des_cipher_top_tb;

architecture behavior of des_cipher_top_tb is

    --=============================================================================================
    -- Constants
    --=============================================================================================
    -- clock period
    constant CLOCK_PERIOD : time := CLK_PERIOD;          -- clock

    --=============================================================================================
    -- Signals
    --=============================================================================================
    --- clock and reset signals ---
    signal clock            : std_logic := '1';                 -- 100MHz clock
    signal reset            : std_logic := '1';                 -- reset active high
    --- input data ---
    signal key_in           : std_logic_vector (0 to 63);   -- key input
    signal data_in          : std_logic_vector (0 to 63);   -- data input
    --- control signals ---
    signal funct_select     : std_logic;                        -- function select: '1' = encryption, '0' = decryption
    signal lddata           : std_logic;                        -- data strobe (active high)
    signal core_busy        : std_logic;
    signal des_out_rdy      : std_logic;
    --- output data ---
    signal data_out         : std_logic_vector (0 to 63);   -- data output

begin

    --=============================================================================================
    -- INSTANTIATION FOR THE DEVICE UNDER TEST
    --=============================================================================================
	Inst_des_cipher_top_dut: entity work.des_cipher_top
        port map(
            --
            -- Core Interface
            --
            key_in            => key_in,            -- input for key

            function_select   => funct_select,      -- function	select: '1' = encryption, '0' = decryption

            data_in           => data_in,           -- input for data

            data_out          => data_out,          -- output for data

            lddata            => lddata,            -- data strobe (active high)
            core_busy         => core_busy,         -- active high when encrypting/decryption data
            des_out_rdy       => des_out_rdy,       -- active high when encryption/decryption of data is done

            reset             => reset,             -- active high
            clock             => clock              -- master clock

        );

    --=============================================================================================
    -- CLOCK GENERATION
    --=============================================================================================
    clock_proc: process is
    begin
        loop
            clock <= not clock;
            wait for CLOCK_PERIOD / 2;
        end loop;
    end process clock_proc;
    --=============================================================================================
    -- TEST BENCH STIMULI
    --=============================================================================================
    -- This testbench exercises the DES toplevel with the 2 test vectors.
    --
    tb1 : process is
    begin
        reset <= '1';
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"6163746976697479";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6d9119c669310aec" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"6d9119c669310aec";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6163746976697479" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"6a617a7a69657374";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"eeea69156ff89f02" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"eeea69156ff89f02";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6a617a7a69657374" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"62757a7a776f7264";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"9c137625bdaf9e2a" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"9c137625bdaf9e2a";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"62757a7a776f7264" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"537461726275636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"2ea7641b231e2879" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"2ea7641b231e2879";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"537461726275636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"666c61706a61636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"fe5999073209146a" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"fe5999073209146a";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"666c61706a61636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"6b69636b6261636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"d2bb0344aa0d2934" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"d2bb0344aa0d2934";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6b69636b6261636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"6261636b7061636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"ca16f578a083ad54" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"ca16f578a083ad54";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6261636b7061636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"70697a7a65726961";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"19164857b1ed1eed" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"19164857b1ed1eed";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"70697a7a65726961" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"6a69756a69747375";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"261259ae6709b30b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"261259ae6709b30b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6a69756a69747375" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"717569786f746963";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"267bb4e213e9cb6c" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"626c697a7a617264";
        funct_select      <= '0';
        data_in           <= X"267bb4e213e9cb6c";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"717569786f746963" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"6163746976697479";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"9f829be191927723" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"9f829be191927723";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6163746976697479" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"6a617a7a69657374";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"5f6025ee951ab781" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"5f6025ee951ab781";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6a617a7a69657374" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"62757a7a776f7264";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"5b30967e0a86728d" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"5b30967e0a86728d";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"62757a7a776f7264" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"537461726275636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"68b01c51d3527994" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"68b01c51d3527994";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"537461726275636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"666c61706a61636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"339c207e9a17ae71" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"339c207e9a17ae71";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"666c61706a61636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"6b69636b6261636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"7f84e8bfcdea91f0" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"7f84e8bfcdea91f0";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6b69636b6261636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"6261636b7061636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"550fa57808371e2e" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"550fa57808371e2e";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6261636b7061636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"70697a7a65726961";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"1102411f6bbc097e" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"1102411f6bbc097e";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"70697a7a65726961" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"6a69756a69747375";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"7db631b575febe1e" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"7db631b575febe1e";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6a69756a69747375" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"717569786f746963";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"b7be9bf61cfc366d" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"736b69706a61636b";
        funct_select      <= '0';
        data_in           <= X"b7be9bf61cfc366d";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"717569786f746963" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"6163746976697479";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"99f8be595bf2f01d" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"99f8be595bf2f01d";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6163746976697479" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"6a617a7a69657374";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"e681d63eba09fe79" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"e681d63eba09fe79";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6a617a7a69657374" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"62757a7a776f7264";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"319b05b610c975ba" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"319b05b610c975ba";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"62757a7a776f7264" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"537461726275636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"74fd27396930e6da" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"74fd27396930e6da";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"537461726275636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"666c61706a61636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"e41718aac3dbf70c" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"e41718aac3dbf70c";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"666c61706a61636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"6b69636b6261636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"e2a8133d7aa58469" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"e2a8133d7aa58469";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6b69636b6261636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"6261636b7061636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"842d91012158c927" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"842d91012158c927";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6261636b7061636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"70697a7a65726961";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"90b3d89867a05f32" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"90b3d89867a05f32";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"70697a7a65726961" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"6a69756a69747375";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"980f94a7e3d89ffe" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"980f94a7e3d89ffe";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6a69756a69747375" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"717569786f746963";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"f6bbaefb29ead11a" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6a756d706f666673";
        funct_select      <= '0';
        data_in           <= X"f6bbaefb29ead11a";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"717569786f746963" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"6163746976697479";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"3a830584d27ad91d" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"3a830584d27ad91d";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6163746976697479" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"6a617a7a69657374";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"bda4bad4688b7560" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"bda4bad4688b7560";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6a617a7a69657374" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"62757a7a776f7264";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"f095bb0f072faec2" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"f095bb0f072faec2";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"62757a7a776f7264" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"537461726275636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"ee92bbaac381752e" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"ee92bbaac381752e";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"537461726275636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"666c61706a61636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"2ca582e5976851e5" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"2ca582e5976851e5";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"666c61706a61636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"6b69636b6261636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"aa9160e33bba4153" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"aa9160e33bba4153";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6b69636b6261636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"6261636b7061636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"bfde88762be7ac83" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"bfde88762be7ac83";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6261636b7061636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"70697a7a65726961";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"b8d57097775af2f2" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"b8d57097775af2f2";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"70697a7a65726961" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"6a69756a69747375";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"f0de212985fe3ec7" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"f0de212985fe3ec7";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6a69756a69747375" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"717569786f746963";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"0a06cbcaae9cf2e9" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"6d6178696d697a65";
        funct_select      <= '0';
        data_in           <= X"0a06cbcaae9cf2e9";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"717569786f746963" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"6163746976697479";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"dee462ec78822bf4" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"dee462ec78822bf4";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6163746976697479" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"6a617a7a69657374";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"118603a096dccc0f" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"118603a096dccc0f";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6a617a7a69657374" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"62757a7a776f7264";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"7858422ded63415c" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"7858422ded63415c";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"62757a7a776f7264" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"537461726275636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"674186b927fd587d" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"674186b927fd587d";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"537461726275636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"666c61706a61636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"57ae29716c76c2ba" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"57ae29716c76c2ba";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"666c61706a61636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"6b69636b6261636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"ae16de56b15e74ef" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"ae16de56b15e74ef";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6b69636b6261636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"6261636b7061636b";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"41fa01ff9afe67e9" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"41fa01ff9afe67e9";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6261636b7061636b" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"70697a7a65726961";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"73ab1ac68adecd0c" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"73ab1ac68adecd0c";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"70697a7a65726961" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"6a69756a69747375";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"48f3065d79a08617" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"48f3065d79a08617";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"6a69756a69747375" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"717569786f746963";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"cb850fb284cb4a9c" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        wait for CLOCK_PERIOD*5;
        reset <= '1';
        wait for CLOCK_PERIOD;
        reset <= '0';
        key_in            <= X"656e67696e656572";
        funct_select      <= '0';
        data_in           <= X"cb850fb284cb4a9c";
        lddata            <= '1';
        wait until des_out_rdy = '1';

        assert data_out = X"717569786f746963" report "test #2 failed" severity error;

        -------------------------------------------------------------------------------------------
        reset <= '1';
                wait; -- stop simulation
            end process tb1;
            --  End Test Bench
        END;
